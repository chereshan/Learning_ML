"row_id","target"
37518,18
37519,18
37520,15
37521,15
37522,18
37523,1
37524,18
37525,18
37526,15
37527,15
37528,18
37529,1
37530,1
37531,1
37532,1
37533,1
37534,3
37535,3
37536,1
37537,1
37538,1
37539,1
37540,1
37541,1
37542,1
37543,1
37544,1
37545,3
37546,3
37547,3
37548,33
37549,33
37550,37
37551,33
37552,33
37553,37
37554,11
37555,33
37556,33
37557,37
37558,11
37559,12
37560,12
37561,11
37562,11
37563,12
37564,11
37565,11
37566,12
37567,12
37568,11
37569,11
37570,37
37571,11
37572,33
37573,33
37574,37
37575,11
37576,11
37577,37
37578,12
37579,49
37580,49
37581,49
37582,49
37583,49
37584,49
37585,49
37586,12
37587,49
37588,49
37589,48
37590,53
37591,53
37592,49
37593,48
37594,53
37595,53
37596,49
37597,53
37598,53
37599,49
37600,48
37601,53
37602,53
37603,49
37604,12
37605,15
37606,15
37607,19
37608,19
37609,15
37610,15
37611,37
37612,12
37613,12
37614,15
37615,15
37616,15
37617,15
37618,15
37619,15
37620,15
37621,37
37622,12
37623,12
37624,12
37625,37
37626,33
37627,33
37628,12
37629,12
37630,12
37631,12
37632,12
37633,12
37634,12
37635,12
37636,33
37637,33
37638,33
37639,33
37640,37
37641,18
37642,18
37643,53
37644,53
37645,37
37646,18
37647,18
37648,9
37649,12
37650,12
37651,37
37652,47
37653,53
37654,53
37655,37
37656,9
37657,12
37658,12
37659,15
37660,19
37661,19
37662,12
37663,12
37664,12
37665,12
37666,19
37667,12
37668,12
37669,53
37670,15
37671,53
37672,15
37673,12
37674,12
37675,12
37676,12
37677,12
37678,15
37679,15
37680,37
37681,12
37682,12
37683,12
37684,18
37685,18
37686,37
37687,12
37688,15
37689,15
37690,15
37691,15
37692,15
37693,49
37694,3
37695,3
37696,3
37697,3
37698,3
37699,3
37700,3
37701,3
37702,3
37703,3
37704,3
37705,3
37706,3
37707,37
37708,3
37709,11
37710,11
37711,47
37712,11
37713,11
37714,47
37715,11
37716,11
37717,49
37718,49
37719,47
37720,11
37721,11
37722,47
37723,11
37724,11
37725,49
37726,49
37727,27
37728,47
37729,11
37730,11
37731,49
37732,48
37733,48
37734,27
37735,33
37736,33
37737,37
37738,49
37739,48
37740,48
37741,49
37742,49
37743,27
37744,27
37745,37
37746,37
37747,37
37748,27
37749,49
37750,33
37751,33
37752,49
37753,49
37754,49
37755,33
37756,33
37757,49
37758,49
37759,33
37760,48
37761,48
37762,27
37763,27
37764,15
37765,3
37766,3
37767,15
37768,15
37769,18
37770,15
37771,3
37772,3
37773,15
37774,1
37775,1
37776,1
37777,1
37778,55
37779,55
37780,1
37781,1
37782,1
37783,1
37784,1
37785,1
37786,1
37787,1
37788,1
37789,1
37790,1
37791,1
37792,1
37793,1
37794,55
37795,55
37796,1
37797,55
37798,55
37799,3
37800,11
37801,33
37802,33
37803,37
37804,12
37805,12
37806,11
37807,11
37808,37
37809,11
37810,33
37811,33
37812,33
37813,33
37814,37
37815,12
37816,12
37817,12
37818,53
37819,49
37820,49
37821,53
37822,53
37823,49
37824,49
37825,49
37826,49
37827,49
37828,49
37829,49
37830,49
37831,53
37832,53
37833,49
37834,48
37835,53
37836,53
37837,49
37838,48
37839,53
37840,53
37841,49
37842,6
37843,6
37844,12
37845,49
37846,49
37847,12
37848,15
37849,15
37850,15
37851,15
37852,19
37853,37
37854,55
37855,55
37856,37
37857,12
37858,12
37859,15
37860,15
37861,37
37862,19
37863,12
37864,12
37865,15
37866,15
37867,37
37868,55
37869,55
37870,37
37871,12
37872,12
37873,12
37874,12
37875,12
37876,12
37877,12
37878,12
37879,12
37880,37
37881,55
37882,55
37883,37
37884,12
37885,55
37886,12
37887,55
37888,12
37889,37
37890,55
37891,55
37892,37
37893,47
37894,33
37895,33
37896,37
37897,47
37898,33
37899,33
37900,47
37901,37
37902,49
37903,49
37904,37
37905,9
37906,12
37907,12
37908,37
37909,12
37910,12
37911,12
37912,12
37913,12
37914,12
37915,12
37916,15
37917,55
37918,55
37919,12
37920,12
37921,12
37922,12
37923,15
37924,55
37925,55
37926,12
37927,12
37928,15
37929,15
37930,15
37931,37
37932,55
37933,55
37934,55
37935,55
37936,37
37937,12
37938,15
37939,15
37940,12
37941,15
37942,15
37943,55
37944,55
37945,12
37946,15
37947,15
37948,55
37949,55
37950,37
37951,12
37952,15
37953,15
37954,15
37955,53
37956,53
37957,37
37958,15
37959,15
37960,15
37961,3
37962,3
37963,3
37964,3
37965,11
37966,11
37967,49
37968,3
37969,37
37970,11
37971,11
37972,3
37973,11
37974,11
37975,3
37976,49
37977,11
37978,11
37979,12
37980,12
37981,37
37982,55
37983,55
37984,37
37985,15
37986,11
37987,11
37988,37
37989,32
37990,32
37991,27
37992,47
37993,11
37994,11
37995,47
37996,11
37997,11
37998,47
37999,11
38000,11
38001,19
38002,19
38003,27
38004,33
38005,48
38006,48
38007,49
38008,49
38009,49
38010,33
38011,48
38012,48
38013,33
38014,48
38015,48
38016,33
38017,27
38018,27
38019,27
38020,33
38021,33
38022,27
38023,27
38024,15
38025,18
38026,18
38027,15
38028,15
38029,18
38030,55
38031,55
38032,1
38033,1
38034,1
38035,1
38036,1
38037,3
38038,55
38039,55
38040,1
38041,1
38042,55
38043,55
38044,3
38045,11
38046,11
38047,37
38048,11
38049,33
38050,33
38051,37
38052,11
38053,12
38054,12
38055,12
38056,11
38057,11
38058,11
38059,37
38060,33
38061,33
38062,37
38063,55
38064,55
38065,37
38066,50
38067,49
38068,49
38069,50
38070,49
38071,53
38072,53
38073,49
38074,53
38075,49
38076,49
38077,49
38078,49
38079,12
38080,49
38081,12
38082,12
38083,12
38084,12
38085,12
38086,53
38087,53
38088,53
38089,49
38090,53
38091,49
38092,49
38093,49
38094,49
38095,49
38096,12
38097,15
38098,15
38099,19
38100,55
38101,55
38102,37
38103,12
38104,15
38105,15
38106,19
38107,55
38108,55
38109,37
38110,33
38111,55
38112,55
38113,37
38114,9
38115,12
38116,12
38117,9
38118,55
38119,55
38120,37
38121,37
38122,12
38123,12
38124,12
38125,15
38126,53
38127,53
38128,12
38129,12
38130,12
38131,12
38132,12
38133,12
38134,12
38135,15
38136,15
38137,37
38138,37
38139,12
38140,15
38141,15
38142,12
38143,15
38144,15
38145,15
38146,55
38147,55
38148,12
38149,15
38150,15
38151,37
38152,3
38153,11
38154,11
38155,3
38156,37
38157,3
38158,11
38159,11
38160,3
38161,11
38162,11
38163,49
38164,3
38165,11
38166,11
38167,55
38168,55
38169,37
38170,37
38171,55
38172,55
38173,37
38174,55
38175,11
38176,11
38177,6
38178,6
38179,37
38180,47
38181,11
38182,11
38183,47
38184,11
38185,11
38186,47
38187,11
38188,11
38189,6
38190,6
38191,27
38192,27
38193,47
38194,11
38195,11
38196,47
38197,11
38198,11
38199,27
38200,27
38201,27
38202,27
38203,27
38204,47
38205,47
38206,47
38207,47
38208,47
38209,15
38210,1
38211,1
38212,15
38213,15
38214,15
38215,1
38216,34
38217,34
38218,1
38219,1
38220,1
38221,1
38222,1
38223,3
38224,1
38225,55
38226,55
38227,1
38228,1
38229,3
38230,26
38231,33
38232,33
38233,37
38234,55
38235,55
38236,37
38237,11
38238,55
38239,55
38240,37
38241,12
38242,11
38243,11
38244,11
38245,12
38246,12
38247,11
38248,11
38249,11
38250,37
38251,11
38252,37
38253,48
38254,48
38255,48
38256,12
38257,48
38258,48
38259,48
38260,12
38261,12
38262,12
38263,12
38264,12
38265,12
38266,12
38267,12
38268,49
38269,49
38270,49
38271,49
38272,12
38273,48
38274,48
38275,48
38276,48
38277,49
38278,49
38279,12
38280,48
38281,48
38282,48
38283,12
38284,48
38285,48
38286,48
38287,12
38288,12
38289,12
38290,12
38291,48
38292,48
38293,48
38294,12
38295,19
38296,55
38297,12
38298,12
38299,12
38300,12
38301,12
38302,12
38303,12
38304,12
38305,19
38306,55
38307,55
38308,12
38309,12
38310,12
38311,12
38312,19
38313,19
38314,19
38315,37
38316,33
38317,55
38318,55
38319,37
38320,12
38321,12
38322,12
38323,12
38324,37
38325,33
38326,12
38327,12
38328,12
38329,12
38330,37
38331,12
38332,12
38333,12
38334,12
38335,55
38336,55
38337,12
38338,12
38339,55
38340,12
38341,55
38342,12
38343,55
38344,12
38345,55
38346,12
38347,37
38348,12
38349,12
38350,12
38351,48
38352,55
38353,55
38354,55
38355,12
38356,12
38357,55
38358,37
38359,12
38360,12
38361,12
38362,48
38363,55
38364,55
38365,12
38366,12
38367,37
38368,37
38369,12
38370,12
38371,12
38372,12
38373,55
38374,55
38375,12
38376,12
38377,12
38378,12
38379,12
38380,55
38381,55
38382,12
38383,12
38384,12
38385,12
38386,19
38387,19
38388,19
38389,12
38390,19
38391,19
38392,19
38393,12
38394,12
38395,12
38396,12
38397,12
38398,12
38399,55
38400,12
38401,12
38402,12
38403,12
38404,12
38405,12
38406,24
38407,12
38408,12
38409,12
38410,12
38411,12
38412,12
38413,12
38414,14
38415,55
38416,55
38417,37
38418,12
38419,12
38420,12
38421,12
38422,12
38423,12
38424,12
38425,12
38426,12
38427,37
38428,3
38429,3
38430,3
38431,3
38432,11
38433,11
38434,3
38435,11
38436,11
38437,3
38438,11
38439,11
38440,26
38441,3
38442,11
38443,11
38444,55
38445,11
38446,11
38447,19
38448,11
38449,55
38450,55
38451,11
38452,19
38453,11
38454,11
38455,19
38456,55
38457,55
38458,27
38459,27
38460,19
38461,11
38462,11
38463,27
38464,27
38465,19
38466,11
38467,11
38468,11
38469,11
38470,27
38471,27
38472,19
38473,11
38474,11
38475,27
38476,37
38477,37
38478,27
38479,48
38480,33
38481,33
38482,27
38483,27
38484,47
38485,49
38486,49
38487,47
38488,47
38489,47
38490,18
38491,18
38492,47
38493,29
38494,29
38495,49
38496,49
38497,15
38498,3
38499,3
38500,15
38501,15
38502,18
38503,3
38504,55
38505,55
38506,1
38507,3
38508,1
38509,1
38510,1
38511,3
38512,55
38513,55
38514,55
38515,11
38516,55
38517,55
38518,37
38519,11
38520,12
38521,12
38522,11
38523,11
38524,37
38525,11
38526,12
38527,11
38528,11
38529,12
38530,12
38531,11
38532,55
38533,11
38534,55
38535,37
38536,12
38537,11
38538,11
38539,12
38540,12
38541,11
38542,11
38543,37
38544,11
38545,12
38546,12
38547,11
38548,11
38549,37
38550,11
38551,55
38552,53
38553,12
38554,32
38555,53
38556,53
38557,12
38558,49
38559,53
38560,53
38561,12
38562,32
38563,32
38564,53
38565,53
38566,12
38567,53
38568,53
38569,12
38570,53
38571,53
38572,12
38573,53
38574,53
38575,53
38576,12
38577,53
38578,53
38579,53
38580,9
38581,19
38582,19
38583,12
38584,12
38585,12
38586,12
38587,12
38588,12
38589,19
38590,19
38591,19
38592,55
38593,55
38594,19
38595,37
38596,55
38597,55
38598,37
38599,12
38600,12
38601,15
38602,15
38603,37
38604,55
38605,55
38606,55
38607,55
38608,55
38609,33
38610,37
38611,37
38612,37
38613,55
38614,55
38615,55
38616,55
38617,55
38618,55
38619,55
38620,55
38621,55
38622,55
38623,37
38624,55
38625,55
38626,55
38627,33
38628,55
38629,55
38630,37
38631,9
38632,33
38633,12
38634,12
38635,9
38636,9
38637,37
38638,9
38639,9
38640,9
38641,37
38642,9
38643,12
38644,12
38645,9
38646,55
38647,55
38648,37
38649,9
38650,55
38651,55
38652,37
38653,9
38654,9
38655,9
38656,32
38657,55
38658,55
38659,12
38660,32
38661,55
38662,55
38663,12
38664,9
38665,55
38666,15
38667,15
38668,37
38669,55
38670,55
38671,55
38672,37
38673,37
38674,12
38675,15
38676,15
38677,12
38678,15
38679,15
38680,14
38681,12
38682,12
38683,15
38684,15
38685,15
38686,15
38687,37
38688,37
38689,9
38690,15
38691,15
38692,3
38693,3
38694,3
38695,3
38696,3
38697,3
38698,3
38699,11
38700,11
38701,55
38702,55
38703,11
38704,55
38705,11
38706,55
38707,11
38708,11
38709,37
38710,55
38711,37
38712,55
38713,37
38714,37
38715,55
38716,11
38717,11
38718,55
38719,11
38720,11
38721,47
38722,11
38723,11
38724,47
38725,11
38726,11
38727,47
38728,11
38729,11
38730,47
38731,11
38732,11
38733,27
38734,27
38735,37
38736,47
38737,11
38738,11
38739,47
38740,11
38741,11
38742,47
38743,11
38744,11
38745,49
38746,47
38747,11
38748,11
38749,27
38750,27
38751,33
38752,29
38753,29
38754,33
38755,29
38756,29
38757,49
38758,49
38759,33
38760,33
38761,29
38762,29
38763,33
38764,49
38765,49
38766,29
38767,29
38768,29
38769,33
38770,32
38771,33
38772,32
38773,33
38774,27
38775,27
38776,15
38777,15
38778,15
38779,15
38780,15
38781,15
38782,3
38783,3
38784,18
38785,15
38786,18
38787,18
38788,15
38789,15
38790,18
38791,3
38792,3
38793,3
38794,11
38795,11
38796,11
38797,37
38798,12
38799,11
38800,11
38801,12
38802,12
38803,11
38804,11
38805,37
38806,11
38807,12
38808,12
38809,11
38810,11
38811,37
38812,11
38813,33
38814,33
38815,37
38816,11
38817,33
38818,33
38819,37
38820,12
38821,0
38822,0
38823,12
38824,12
38825,11
38826,11
38827,37
38828,11
38829,33
38830,33
38831,33
38832,37
38833,11
38834,12
38835,12
38836,11
38837,11
38838,37
38839,11
38840,11
38841,11
38842,11
38843,11
38844,37
38845,32
38846,49
38847,49
38848,49
38849,32
38850,53
38851,53
38852,49
38853,32
38854,49
38855,53
38856,53
38857,49
38858,49
38859,49
38860,49
38861,49
38862,53
38863,53
38864,53
38865,49
38866,12
38867,12
38868,12
38869,48
38870,49
38871,49
38872,53
38873,53
38874,49
38875,49
38876,12
38877,19
38878,12
38879,12
38880,15
38881,15
38882,37
38883,12
38884,15
38885,15
38886,19
38887,19
38888,19
38889,19
38890,37
38891,12
38892,33
38893,33
38894,12
38895,12
38896,12
38897,33
38898,33
38899,37
38900,9
38901,12
38902,12
38903,49
38904,49
38905,37
38906,9
38907,12
38908,0
38909,12
38910,0
38911,53
38912,53
38913,53
38914,53
38915,37
38916,47
38917,53
38918,53
38919,37
38920,15
38921,15
38922,19
38923,19
38924,15
38925,12
38926,12
38927,12
38928,12
38929,12
38930,12
38931,12
38932,15
38933,15
38934,12
38935,12
38936,12
38937,12
38938,12
38939,12
38940,15
38941,15
38942,12
38943,12
38944,12
38945,12
38946,12
38947,12
38948,12
38949,15
38950,15
38951,15
38952,37
38953,12
38954,12
38955,12
38956,15
38957,15
38958,15
38959,12
38960,12
38961,53
38962,53
38963,15
38964,15
38965,37
38966,37
38967,37
38968,37
38969,3
38970,3
38971,0
38972,3
38973,0
38974,15
38975,15
38976,37
38977,3
38978,3
38979,3
38980,3
38981,3
38982,3
38983,3
38984,3
38985,0
38986,3
38987,0
38988,3
38989,3
38990,3
38991,3
38992,3
38993,3
38994,3
38995,3
38996,3
38997,3
38998,3
38999,3
39000,3
39001,3
39002,3
39003,47
39004,11
39005,11
39006,49
39007,49
39008,47
39009,11
39010,11
39011,47
39012,11
39013,11
39014,47
39015,11
39016,11
39017,33
39018,33
39019,33
39020,49
39021,49
39022,29
39023,48
39024,48
39025,37
39026,37
39027,33
39028,48
39029,48
39030,27
39031,27
39032,27
39033,33
39034,33
39035,33
39036,33
39037,27
39038,27
39039,48
39040,48
39041,47
39042,47
39043,47
39044,47
39045,47
39046,15
39047,3
39048,3
39049,15
39050,15
39051,15
39052,15
39053,3
39054,3
39055,15
39056,3
39057,1
39058,1
39059,1
39060,3
39061,1
39062,1
39063,1
39064,1
39065,3
39066,3
39067,55
39068,55
39069,3
39070,11
39071,12
39072,12
39073,11
39074,11
39075,37
39076,11
39077,33
39078,33
39079,37
39080,11
39081,12
39082,12
39083,11
39084,11
39085,37
39086,11
39087,12
39088,12
39089,11
39090,11
39091,37
39092,12
39093,11
39094,11
39095,12
39096,12
39097,11
39098,11
39099,37
39100,49
39101,33
39102,33
39103,37
39104,37
39105,37
39106,37
39107,53
39108,53
39109,12
39110,53
39111,53
39112,12
39113,53
39114,53
39115,48
39116,53
39117,53
39118,49
39119,53
39120,53
39121,49
39122,49
39123,49
39124,12
39125,12
39126,12
39127,48
39128,53
39129,53
39130,49
39131,48
39132,53
39133,53
39134,49
39135,19
39136,12
39137,12
39138,15
39139,15
39140,37
39141,12
39142,15
39143,15
39144,55
39145,55
39146,37
39147,12
39148,12
39149,33
39150,55
39151,55
39152,37
39153,12
39154,12
39155,12
39156,55
39157,55
39158,33
39159,9
39160,12
39161,12
39162,49
39163,49
39164,15
39165,15
39166,37
39167,47
39168,47
39169,15
39170,15
39171,55
39172,55
39173,37
39174,55
39175,55
39176,37
39177,9
39178,55
39179,55
39180,47
39181,49
39182,49
39183,37
39184,15
39185,53
39186,53
39187,12
39188,12
39189,12
39190,12
39191,12
39192,12
39193,12
39194,55
39195,55
39196,12
39197,12
39198,12
39199,19
39200,53
39201,53
39202,12
39203,15
39204,55
39205,15
39206,15
39207,55
39208,15
39209,12
39210,55
39211,55
39212,12
39213,55
39214,15
39215,15
39216,55
39217,37
39218,55
39219,55
39220,37
39221,15
39222,15
39223,15
39224,15
39225,15
39226,15
39227,15
39228,55
39229,55
39230,37
39231,37
39232,37
39233,15
39234,15
39235,15
39236,3
39237,3
39238,3
39239,3
39240,3
39241,3
39242,15
39243,15
39244,37
39245,3
39246,3
39247,3
39248,3
39249,3
39250,3
39251,3
39252,3
39253,11
39254,11
39255,3
39256,11
39257,11
39258,6
39259,6
39260,3
39261,11
39262,11
39263,55
39264,11
39265,11
39266,55
39267,11
39268,11
39269,47
39270,11
39271,11
39272,49
39273,47
39274,11
39275,11
39276,11
39277,11
39278,47
39279,11
39280,11
39281,19
39282,19
39283,27
39284,47
39285,11
39286,11
39287,47
39288,6
39289,6
39290,47
39291,11
39292,11
39293,47
39294,11
39295,11
39296,47
39297,27
39298,27
39299,27
39300,27
39301,27
39302,27
39303,27
39304,47
39305,11
39306,11
39307,33
39308,29
39309,29
39310,37
39311,37
39312,27
39313,48
39314,48
39315,48
39316,27
39317,27
39318,48
39319,48
39320,48
39321,33
39322,33
39323,33
39324,27
39325,27
39326,15
39327,15
39328,15
39329,15
39330,15
39331,15
39332,15
39333,15
39334,15
39335,15
39336,15
39337,15
39338,15
39339,15
39340,3
39341,18
39342,18
39343,15
39344,15
39345,18
39346,15
39347,3
39348,3
39349,18
39350,1
39351,1
39352,1
39353,1
39354,3
39355,1
39356,1
39357,3
39358,3
39359,33
39360,33
39361,37
39362,11
39363,12
39364,12
39365,11
39366,11
39367,37
39368,11
39369,11
39370,55
39371,55
39372,11
39373,37
39374,12
39375,55
39376,55
39377,12
39378,12
39379,11
39380,11
39381,37
39382,32
39383,49
39384,49
39385,49
39386,49
39387,12
39388,49
39389,53
39390,53
39391,12
39392,12
39393,53
39394,53
39395,12
39396,12
39397,12
39398,49
39399,49
39400,49
39401,49
39402,12
39403,50
39404,49
39405,49
39406,12
39407,50
39408,49
39409,49
39410,12
39411,50
39412,53
39413,53
39414,12
39415,50
39416,53
39417,53
39418,12
39419,50
39420,6
39421,6
39422,53
39423,53
39424,12
39425,19
39426,19
39427,53
39428,49
39429,49
39430,49
39431,49
39432,49
39433,49
39434,37
39435,53
39436,53
39437,53
39438,37
39439,12
39440,15
39441,15
39442,19
39443,55
39444,55
39445,37
39446,15
39447,15
39448,12
39449,19
39450,15
39451,15
39452,55
39453,55
39454,37
39455,19
39456,54
39457,54
39458,15
39459,15
39460,37
39461,33
39462,55
39463,55
39464,37
39465,55
39466,55
39467,55
39468,55
39469,55
39470,55
39471,33
39472,55
39473,55
39474,37
39475,9
39476,12
39477,12
39478,9
39479,12
39480,12
39481,37
39482,33
39483,15
39484,15
39485,37
39486,9
39487,12
39488,12
39489,9
39490,9
39491,37
39492,9
39493,12
39494,55
39495,12
39496,55
39497,9
39498,9
39499,9
39500,37
39501,37
39502,12
39503,12
39504,12
39505,15
39506,15
39507,55
39508,55
39509,12
39510,15
39511,55
39512,15
39513,55
39514,12
39515,12
39516,12
39517,12
39518,55
39519,55
39520,55
39521,12
39522,37
39523,12
39524,12
39525,55
39526,55
39527,55
39528,37
39529,55
39530,15
39531,15
39532,37
39533,55
39534,15
39535,15
39536,37
39537,37
39538,15
39539,15
39540,15
39541,14
39542,55
39543,55
39544,37
39545,15
39546,15
39547,15
39548,15
39549,15
39550,15
39551,37
39552,37
39553,37
39554,15
39555,15
39556,15
39557,37
39558,37
39559,3
39560,3
39561,3
39562,3
39563,3
39564,3
39565,55
39566,37
39567,3
39568,3
39569,3
39570,3
39571,3
39572,3
39573,3
39574,11
39575,11
39576,19
39577,19
39578,3
39579,11
39580,55
39581,55
39582,11
39583,3
39584,11
39585,11
39586,55
39587,11
39588,11
39589,55
39590,11
39591,55
39592,11
39593,55
39594,6
39595,6
39596,47
39597,11
39598,11
39599,19
39600,11
39601,11
39602,27
39603,27
39604,19
39605,19
39606,11
39607,11
39608,27
39609,27
39610,11
39611,11
39612,49
39613,29
39614,29
39615,29
39616,54
39617,54
39618,29
39619,29
39620,29
39621,33
39622,33
39623,27
39624,27
39625,29
39626,29
39627,33
39628,29
39629,33
39630,29
39631,29
39632,33
39633,27
39634,33
39635,27
39636,33
39637,27
39638,27
39639,29
39640,29
39641,29
39642,33
39643,33
39644,27
39645,27
39646,29
39647,29
39648,33
39649,29
39650,33
39651,27
39652,27
39653,18
39654,18
39655,18
39656,18
39657,18
39658,3
39659,1
39660,1
39661,3
39662,1
39663,55
39664,55
39665,3
39666,3
39667,1
39668,1
39669,3
39670,1
39671,3
39672,3
39673,3
39674,3
39675,1
39676,1
39677,3
39678,3
39679,1
39680,1
39681,3
39682,33
39683,33
39684,33
39685,37
39686,33
39687,33
39688,37
39689,11
39690,11
39691,37
39692,26
39693,12
39694,12
39695,11
39696,11
39697,37
39698,11
39699,32
39700,32
39701,12
39702,12
39703,12
39704,12
39705,12
39706,12
39707,12
39708,12
39709,12
39710,48
39711,53
39712,53
39713,12
39714,48
39715,12
39716,12
39717,12
39718,53
39719,53
39720,12
39721,48
39722,53
39723,53
39724,12
39725,48
39726,12
39727,12
39728,24
39729,24
39730,53
39731,12
39732,53
39733,12
39734,12
39735,12
39736,12
39737,12
39738,12
39739,12
39740,12
39741,12
39742,12
39743,12
39744,12
39745,12
39746,48
39747,48
39748,48
39749,12
39750,12
39751,12
39752,12
39753,12
39754,12
39755,55
39756,12
39757,55
39758,55
39759,55
39760,12
39761,19
39762,55
39763,55
39764,12
39765,55
39766,55
39767,12
39768,12
39769,18
39770,18
39771,12
39772,12
39773,12
39774,12
39775,12
39776,12
39777,37
39778,19
39779,55
39780,55
39781,37
39782,19
39783,19
39784,12
39785,12
39786,12
39787,55
39788,37
39789,37
39790,19
39791,19
39792,19
39793,37
39794,12
39795,12
39796,12
39797,55
39798,37
39799,37
39800,37
39801,12
39802,12
39803,12
39804,33
39805,12
39806,12
39807,37
39808,12
39809,12
39810,12
39811,33
39812,55
39813,55
39814,37
39815,48
39816,12
39817,12
39818,37
39819,19
39820,19
39821,12
39822,12
39823,12
39824,12
39825,12
39826,12
39827,12
39828,12
39829,12
39830,12
39831,19
39832,55
39833,55
39834,12
39835,19
39836,19
39837,19
39838,12
39839,19
39840,19
39841,19
39842,12
39843,19
39844,19
39845,19
39846,12
39847,12
39848,55
39849,55
39850,55
39851,12
39852,12
39853,12
39854,12
39855,12
39856,12
39857,12
39858,12
39859,12
39860,12
39861,12
39862,55
39863,12
39864,55
39865,12
39866,12
39867,12
39868,12
39869,12
39870,12
39871,12
39872,12
39873,12
39874,12
39875,24
39876,55
39877,55
39878,55
39879,12
39880,12
39881,12
39882,12
39883,12
39884,55
39885,55
39886,12
39887,12
39888,12
39889,12
39890,12
39891,12
39892,12
39893,12
39894,12
39895,12
39896,12
39897,12
39898,12
39899,12
39900,12
39901,55
39902,12
39903,12
39904,55
39905,55
39906,12
39907,12
39908,12
39909,12
39910,12
39911,55
39912,55
39913,12
39914,12
39915,55
39916,37
39917,37
39918,37
39919,37
39920,3
39921,3
39922,3
39923,12
39924,12
39925,37
39926,37
39927,3
39928,6
39929,6
39930,12
39931,12
39932,3
39933,55
39934,3
39935,55
39936,3
39937,12
39938,12
39939,26
39940,55
39941,3
39942,3
39943,12
39944,12
39945,26
39946,27
39947,27
39948,27
39949,27
39950,27
39951,27
39952,27
39953,27
39954,27
39955,27
39956,27
39957,27
39958,27
39959,27
39960,27
39961,27
39962,27
39963,27
39964,27
39965,27
39966,27
39967,27
39968,27
39969,27
39970,27
39971,27
39972,27
39973,27
39974,33
39975,48
39976,48
39977,27
39978,27
39979,27
39980,27
39981,27
39982,27
39983,27
39984,27
39985,27
39986,27
39987,47
39988,47
39989,47
39990,47
39991,37
39992,37
39993,47
39994,47
39995,47
39996,47
39997,47
39998,47
39999,47
40000,47
40001,1
40002,18
40003,18
40004,49
40005,18
40006,18
40007,1
40008,1
40009,6
40010,1
40011,1
40012,1
40013,1
40014,1
40015,1
40016,1
40017,6
40018,1
40019,6
40020,1
40021,6
40022,6
40023,18
40024,18
40025,1
40026,1
40027,6
40028,1
40029,1
40030,1
40031,6
40032,6
40033,6
40034,6
40035,6
40036,6
40037,37
40038,37
40039,37
40040,47
40041,6
40042,6
40043,49
40044,49
40045,55
40046,12
40047,12
40048,37
40049,37
40050,37
40051,55
40052,19
40053,19
40054,12
40055,12
40056,12
40057,12
40058,12
40059,18
40060,18
40061,15
40062,15
40063,18
40064,3
40065,1
40066,1
40067,1
40068,1
40069,3
40070,1
40071,1
40072,1
40073,1
40074,3
40075,1
40076,1
40077,1
40078,1
40079,3
40080,3
40081,1
40082,1
40083,3
40084,3
40085,3
40086,3
40087,3
40088,3
40089,1
40090,1
40091,3
40092,33
40093,12
40094,11
40095,11
40096,12
40097,12
40098,11
40099,11
40100,33
40101,33
40102,37
40103,33
40104,33
40105,37
40106,11
40107,12
40108,12
40109,11
40110,11
40111,37
40112,11
40113,11
40114,11
40115,37
40116,37
40117,11
40118,11
40119,37
40120,37
40121,12
40122,12
40123,11
40124,11
40125,37
40126,33
40127,33
40128,37
40129,37
40130,33
40131,33
40132,37
40133,12
40134,12
40135,49
40136,49
40137,12
40138,12
40139,12
40140,12
40141,32
40142,53
40143,53
40144,12
40145,32
40146,32
40147,53
40148,53
40149,12
40150,53
40151,53
40152,12
40153,32
40154,53
40155,53
40156,12
40157,32
40158,53
40159,53
40160,12
40161,18
40162,12
40163,12
40164,19
40165,19
40166,19
40167,19
40168,19
40169,37
40170,37
40171,19
40172,12
40173,12
40174,15
40175,15
40176,37
40177,15
40178,15
40179,19
40180,19
40181,19
40182,37
40183,15
40184,15
40185,15
40186,12
40187,12
40188,12
40189,33
40190,12
40191,12
40192,37
40193,33
40194,37
40195,33
40196,37
40197,12
40198,12
40199,12
40200,12
40201,33
40202,33
40203,12
40204,9
40205,12
40206,12
40207,9
40208,12
40209,12
40210,12
40211,12
40212,15
40213,15
40214,37
40215,33
40216,33
40217,37
40218,47
40219,53
40220,15
40221,15
40222,53
40223,53
40224,53
40225,37
40226,15
40227,15
40228,37
40229,9
40230,12
40231,12
40232,47
40233,53
40234,53
40235,49
40236,37
40237,18
40238,18
40239,37
40240,49
40241,15
40242,15
40243,12
40244,19
40245,19
40246,12
40247,12
40248,12
40249,15
40250,15
40251,12
40252,12
40253,12
40254,12
40255,19
40256,19
40257,19
40258,12
40259,12
40260,12
40261,15
40262,15
40263,15
40264,15
40265,15
40266,37
40267,15
40268,37
40269,15
40270,15
40271,15
40272,15
40273,53
40274,53
40275,3
40276,3
40277,3
40278,3
40279,3
40280,3
40281,37
40282,3
40283,0
40284,0
40285,3
40286,3
40287,6
40288,3
40289,6
40290,3
40291,3
40292,3
40293,3
40294,3
40295,3
40296,3
40297,49
40298,3
40299,3
40300,47
40301,11
40302,11
40303,47
40304,47
40305,47
40306,11
40307,11
40308,37
40309,19
40310,19
40311,11
40312,11
40313,11
40314,11
40315,19
40316,11
40317,11
40318,19
40319,11
40320,11
40321,32
40322,29
40323,29
40324,32
40325,29
40326,29
40327,33
40328,33
40329,33
40330,27
40331,27
40332,33
40333,32
40334,32
40335,27
40336,27
40337,33
40338,32
40339,32
40340,33
40341,33
40342,27
40343,27
40344,27
40345,27
40346,27
40347,27
40348,27
40349,27
40350,27
40351,1
40352,55
40353,55
40354,1
40355,1
40356,55
40357,55
40358,1
40359,1
40360,1
40361,1
40362,1
40363,3
40364,1
40365,1
40366,1
40367,3
40368,1
40369,1
40370,1
40371,1
40372,3
40373,33
40374,33
40375,33
40376,37
40377,11
40378,33
40379,33
40380,37
40381,33
40382,33
40383,37
40384,11
40385,12
40386,0
40387,0
40388,12
40389,12
40390,11
40391,11
40392,33
40393,33
40394,37
40395,11
40396,55
40397,55
40398,37
40399,53
40400,53
40401,12
40402,32
40403,49
40404,49
40405,49
40406,49
40407,12
40408,32
40409,53
40410,53
40411,12
40412,32
40413,49
40414,32
40415,49
40416,49
40417,12
40418,53
40419,32
40420,53
40421,12
40422,49
40423,49
40424,53
40425,53
40426,49
40427,49
40428,12
40429,32
40430,49
40431,49
40432,12
40433,12
40434,12
40435,12
40436,32
40437,49
40438,53
40439,53
40440,49
40441,49
40442,12
40443,12
40444,49
40445,49
40446,49
40447,49
40448,12
40449,49
40450,49
40451,53
40452,6
40453,6
40454,19
40455,19
40456,19
40457,19
40458,19
40459,19
40460,12
40461,15
40462,15
40463,19
40464,55
40465,55
40466,37
40467,6
40468,6
40469,55
40470,6
40471,6
40472,19
40473,19
40474,55
40475,55
40476,55
40477,37
40478,55
40479,55
40480,37
40481,37
40482,19
40483,19
40484,55
40485,55
40486,55
40487,55
40488,55
40489,55
40490,55
40491,55
40492,55
40493,55
40494,12
40495,12
40496,0
40497,0
40498,12
40499,12
40500,9
40501,12
40502,12
40503,55
40504,55
40505,37
40506,15
40507,15
40508,55
40509,15
40510,55
40511,15
40512,37
40513,47
40514,55
40515,55
40516,37
40517,9
40518,12
40519,12
40520,47
40521,9
40522,55
40523,15
40524,55
40525,15
40526,55
40527,15
40528,55
40529,12
40530,15
40531,12
40532,37
40533,47
40534,55
40535,55
40536,9
40537,47
40538,55
40539,55
40540,55
40541,55
40542,37
40543,37
40544,37
40545,19
40546,19
40547,19
40548,53
40549,53
40550,12
40551,12
40552,55
40553,12
40554,55
40555,12
40556,55
40557,55
40558,15
40559,15
40560,12
40561,55
40562,55
40563,15
40564,15
40565,55
40566,55
40567,12
40568,12
40569,12
40570,6
40571,6
40572,19
40573,19
40574,55
40575,55
40576,55
40577,55
40578,15
40579,15
40580,19
40581,19
40582,55
40583,19
40584,19
40585,15
40586,15
40587,15
40588,15
40589,15
40590,15
40591,37
40592,37
40593,15
40594,15
40595,15
40596,19
40597,19
40598,3
40599,0
40600,0
40601,3
40602,3
40603,3
40604,1
40605,3
40606,3
40607,3
40608,3
40609,55
40610,3
40611,55
40612,3
40613,55
40614,55
40615,37
40616,55
40617,37
40618,55
40619,37
40620,55
40621,55
40622,37
40623,3
40624,3
40625,3
40626,6
40627,6
40628,55
40629,11
40630,11
40631,55
40632,11
40633,11
40634,55
40635,19
40636,19
40637,11
40638,11
40639,49
40640,47
40641,11
40642,11
40643,19
40644,11
40645,11
40646,19
40647,19
40648,11
40649,11
40650,11
40651,11
40652,19
40653,11
40654,11
40655,19
40656,6
40657,6
40658,19
40659,11
40660,11
40661,11
40662,11
40663,27
40664,27
40665,49
40666,19
40667,11
40668,11
40669,27
40670,27
40671,33
40672,29
40673,29
40674,33
40675,29
40676,33
40677,29
40678,33
40679,27
40680,27
40681,15
40682,15
40683,15
40684,15
40685,15
40686,15
40687,15
40688,18
40689,18
40690,15
40691,15
40692,18
40693,15
40694,3
40695,3
40696,18
40697,1
40698,1
40699,1
40700,1
40701,1
40702,1
40703,3
40704,3
40705,1
40706,1
40707,3
40708,55
40709,55
40710,3
40711,1
40712,33
40713,33
40714,37
40715,33
40716,33
40717,33
40718,33
40719,37
40720,12
40721,12
40722,11
40723,11
40724,37
40725,11
40726,11
40727,37
40728,33
40729,12
40730,12
40731,11
40732,37
40733,12
40734,12
40735,11
40736,11
40737,33
40738,33
40739,11
40740,11
40741,37
40742,11
40743,12
40744,12
40745,11
40746,11
40747,37
40748,11
40749,55
40750,55
40751,37
40752,11
40753,55
40754,55
40755,37
40756,6
40757,6
40758,53
40759,53
40760,53
40761,53
40762,32
40763,53
40764,53
40765,12
40766,12
40767,12
40768,53
40769,49
40770,49
40771,37
40772,53
40773,49
40774,49
40775,49
40776,49
40777,37
40778,18
40779,18
40780,12
40781,15
40782,15
40783,37
40784,19
40785,55
40786,55
40787,37
40788,12
40789,15
40790,15
40791,55
40792,55
40793,37
40794,19
40795,55
40796,55
40797,37
40798,33
40799,55
40800,55
40801,37
40802,37
40803,37
40804,37
40805,55
40806,55
40807,55
40808,55
40809,55
40810,55
40811,55
40812,9
40813,12
40814,12
40815,55
40816,55
40817,37
40818,37
40819,37
40820,55
40821,37
40822,55
40823,55
40824,55
40825,37
40826,37
40827,37
40828,9
40829,9
40830,9
40831,37
40832,37
40833,55
40834,55
40835,37
40836,55
40837,55
40838,37
40839,9
40840,9
40841,9
40842,9
40843,55
40844,9
40845,9
40846,55
40847,9
40848,9
40849,9
40850,32
40851,55
40852,55
40853,12
40854,19
40855,55
40856,55
40857,37
40858,19
40859,19
40860,37
40861,6
40862,6
40863,12
40864,12
40865,12
40866,12
40867,12
40868,12
40869,19
40870,19
40871,15
40872,15
40873,37
40874,19
40875,19
40876,37
40877,37
40878,37
40879,19
40880,19
40881,15
40882,15
40883,55
40884,15
40885,55
40886,55
40887,55
40888,14
40889,14
40890,37
40891,15
40892,15
40893,15
40894,15
40895,15
40896,15
40897,18
40898,18
40899,3
40900,18
40901,18
40902,3
40903,3
40904,3
40905,3
40906,55
40907,55
40908,3
40909,3
40910,3
40911,18
40912,18
40913,3
40914,3
40915,3
40916,18
40917,18
40918,37
40919,3
40920,3
40921,3
40922,55
40923,3
40924,3
40925,3
40926,37
40927,55
40928,55
40929,37
40930,55
40931,3
40932,3
40933,32
40934,11
40935,11
40936,6
40937,6
40938,6
40939,6
40940,27
40941,37
40942,19
40943,11
40944,11
40945,19
40946,49
40947,19
40948,6
40949,6
40950,11
40951,11
40952,19
40953,11
40954,11
40955,33
40956,29
40957,29
40958,33
40959,29
40960,29
40961,29
40962,29
40963,29
40964,54
40965,54
40966,29
40967,29
40968,29
40969,54
40970,54
40971,29
40972,29
40973,29
40974,27
40975,27
40976,27
40977,33
40978,33
40979,27
40980,27
40981,47
40982,47
40983,47
40984,47
40985,47
40986,3
40987,18
40988,18
40989,18
40990,18
40991,18
40992,1
40993,1
40994,1
40995,1
40996,1
40997,1
40998,3
40999,1
41000,1
41001,3
41002,3
41003,55
41004,55
41005,3
41006,3
41007,3
41008,3
41009,1
41010,1
41011,3
41012,1
41013,1
41014,1
41015,1
41016,37
41017,18
41018,18
41019,12
41020,12
41021,11
41022,11
41023,37
41024,12
41025,12
41026,11
41027,11
41028,37
41029,12
41030,55
41031,12
41032,55
41033,12
41034,12
41035,11
41036,11
41037,11
41038,11
41039,37
41040,33
41041,11
41042,11
41043,37
41044,33
41045,12
41046,12
41047,11
41048,11
41049,37
41050,24
41051,55
41052,55
41053,37
41054,33
41055,55
41056,55
41057,37
41058,11
41059,55
41060,55
41061,37
41062,32
41063,32
41064,32
41065,12
41066,32
41067,53
41068,53
41069,12
41070,32
41071,53
41072,53
41073,12
41074,6
41075,6
41076,12
41077,12
41078,48
41079,53
41080,53
41081,12
41082,48
41083,53
41084,53
41085,12
41086,19
41087,12
41088,12
41089,12
41090,12
41091,55
41092,19
41093,12
41094,12
41095,55
41096,19
41097,55
41098,55
41099,37
41100,12
41101,12
41102,12
41103,12
41104,12
41105,37
41106,55
41107,12
41108,12
41109,37
41110,37
41111,37
41112,55
41113,55
41114,55
41115,55
41116,55
41117,55
41118,55
41119,55
41120,55
41121,55
41122,55
41123,55
41124,37
41125,55
41126,37
41127,55
41128,37
41129,18
41130,18
41131,12
41132,12
41133,12
41134,37
41135,33
41136,12
41137,12
41138,55
41139,55
41140,55
41141,55
41142,37
41143,12
41144,12
41145,12
41146,12
41147,12
41148,12
41149,12
41150,12
41151,12
41152,12
41153,12
41154,12
41155,19
41156,55
41157,55
41158,12
41159,19
41160,55
41161,12
41162,55
41163,12
41164,12
41165,12
41166,12
41167,12
41168,12
41169,12
41170,12
41171,12
41172,12
41173,12
41174,12
41175,12
41176,19
41177,12
41178,12
41179,12
41180,19
41181,19
41182,19
41183,19
41184,19
41185,12
41186,19
41187,19
41188,55
41189,55
41190,55
41191,55
41192,12
41193,12
41194,12
41195,55
41196,24
41197,12
41198,12
41199,12
41200,55
41201,12
41202,12
41203,55
41204,12
41205,55
41206,12
41207,12
41208,55
41209,12
41210,55
41211,55
41212,55
41213,55
41214,55
41215,55
41216,55
41217,55
41218,12
41219,12
41220,55
41221,19
41222,19
41223,55
41224,6
41225,6
41226,12
41227,12
41228,12
41229,19
41230,19
41231,12
41232,55
41233,55
41234,12
41235,12
41236,12
41237,12
41238,12
41239,12
41240,12
41241,12
41242,12
41243,3
41244,3
41245,3
41246,18
41247,18
41248,37
41249,3
41250,3
41251,3
41252,3
41253,3
41254,3
41255,37
41256,37
41257,37
41258,3
41259,3
41260,3
41261,55
41262,55
41263,55
41264,55
41265,55
41266,55
41267,19
41268,11
41269,11
41270,19
41271,11
41272,11
41273,19
41274,19
41275,27
41276,19
41277,11
41278,11
41279,27
41280,27
41281,19
41282,11
41283,11
41284,27
41285,27
41286,19
41287,55
41288,55
41289,27
41290,27
41291,33
41292,48
41293,48
41294,26
41295,33
41296,48
41297,48
41298,37
41299,37
41300,27
41301,33
41302,48
41303,48
41304,27
41305,33
41306,27
41307,27
41308,33
41309,27
41310,27
41311,27
41312,27
41313,47
41314,47
41315,37
41316,37
41317,37
41318,37
41319,37
41320,37
41321,47
41322,47
41323,47
41324,47
41325,47
41326,47
41327,47
41328,47
41329,47
41330,47
41331,29
41332,6
41333,6
41334,47
41335,47
41336,6
41337,18
41338,18
41339,6
41340,6
41341,6
41342,6
41343,6
41344,6
41345,6
41346,15
41347,6
41348,6
41349,6
41350,6
41351,19
41352,6
41353,6
41354,15
41355,15
41356,6
41357,19
41358,19
41359,19
41360,19
41361,6
41362,18
41363,18
41364,18
41365,18
41366,19
41367,19
41368,19
41369,19
41370,19
41371,19
41372,15
41373,19
41374,19
41375,6
41376,6
41377,19
41378,19
41379,6
41380,6
41381,18
41382,18
41383,6
41384,6
41385,19
41386,19
41387,47
41388,19
41389,19
41390,49
41391,49
41392,3
41393,1
41394,1
41395,1
41396,1
41397,1
41398,1
41399,1
41400,1
41401,1
41402,1
41403,3
41404,1
41405,3
41406,3
41407,1
41408,1
41409,3
41410,55
41411,55
41412,55
41413,55
41414,55
41415,55
41416,37
41417,33
41418,55
41419,55
41420,37
41421,12
41422,12
41423,11
41424,11
41425,37
41426,37
41427,55
41428,55
41429,37
41430,32
41431,32
41432,32
41433,6
41434,32
41435,32
41436,32
41437,6
41438,32
41439,32
41440,6
41441,32
41442,12
41443,12
41444,6
41445,6
41446,6
41447,32
41448,12
41449,12
41450,12
41451,12
41452,6
41453,19
41454,19
41455,6
41456,6
41457,6
41458,32
41459,53
41460,53
41461,37
41462,12
41463,53
41464,53
41465,55
41466,12
41467,12
41468,15
41469,15
41470,37
41471,55
41472,55
41473,55
41474,37
41475,19
41476,19
41477,18
41478,18
41479,55
41480,55
41481,55
41482,55
41483,55
41484,55
41485,55
41486,37
41487,37
41488,37
41489,18
41490,18
41491,55
41492,55
41493,9
41494,9
41495,37
41496,9
41497,55
41498,55
41499,9
41500,37
41501,9
41502,9
41503,9
41504,9
41505,9
41506,9
41507,55
41508,55
41509,37
41510,32
41511,32
41512,32
41513,12
41514,32
41515,55
41516,55
41517,37
41518,6
41519,6
41520,19
41521,19
41522,55
41523,6
41524,6
41525,15
41526,15
41527,55
41528,55
41529,55
41530,55
41531,55
41532,55
41533,55
41534,55
41535,15
41536,15
41537,55
41538,55
41539,55
41540,55
41541,55
41542,12
41543,15
41544,15
41545,14
41546,14
41547,14
41548,14
41549,37
41550,37
41551,37
41552,19
41553,19
41554,3
41555,3
41556,3
41557,55
41558,3
41559,3
41560,6
41561,6
41562,55
41563,3
41564,3
41565,55
41566,19
41567,19
41568,55
41569,37
41570,37
41571,32
41572,11
41573,55
41574,11
41575,11
41576,55
41577,11
41578,6
41579,6
41580,32
41581,11
41582,11
41583,49
41584,6
41585,6
41586,32
41587,11
41588,11
41589,19
41590,19
41591,6
41592,6
41593,19
41594,19
41595,19
41596,11
41597,11
41598,19
41599,37
41600,37
41601,32
41602,32
41603,32
41604,33
41605,33
41606,32
41607,32
41608,32
41609,33
41610,33
41611,32
41612,32
41613,32
41614,32
41615,29
41616,29
41617,33
41618,33
41619,29
41620,29
41621,29
41622,29
41623,33
41624,33
41625,33
41626,33
41627,33
41628,33
41629,18
41630,18
41631,15
41632,15
41633,18
41634,15
41635,18
41636,18
41637,15
41638,15
41639,18
41640,3
41641,3
41642,3
41643,3
41644,49
41645,12
41646,12
41647,11
41648,11
41649,37
41650,37
41651,11
41652,11
41653,37
41654,37
41655,12
41656,11
41657,11
41658,12
41659,12
41660,11
41661,11
41662,49
41663,37
41664,12
41665,12
41666,11
41667,11
41668,37
41669,12
41670,12
41671,37
41672,37
41673,33
41674,33
41675,37
41676,32
41677,32
41678,32
41679,12
41680,32
41681,32
41682,32
41683,12
41684,32
41685,18
41686,49
41687,18
41688,49
41689,12
41690,32
41691,32
41692,53
41693,53
41694,12
41695,49
41696,49
41697,53
41698,53
41699,49
41700,49
41701,12
41702,32
41703,19
41704,19
41705,53
41706,53
41707,12
41708,32
41709,53
41710,53
41711,12
41712,32
41713,53
41714,53
41715,12
41716,32
41717,49
41718,49
41719,12
41720,6
41721,6
41722,12
41723,12
41724,12
41725,53
41726,53
41727,37
41728,12
41729,12
41730,12
41731,49
41732,49
41733,19
41734,19
41735,37
41736,19
41737,18
41738,18
41739,15
41740,15
41741,37
41742,37
41743,15
41744,15
41745,15
41746,18
41747,18
41748,18
41749,18
41750,12
41751,12
41752,12
41753,9
41754,12
41755,33
41756,12
41757,12
41758,33
41759,12
41760,12
41761,12
41762,47
41763,32
41764,32
41765,37
41766,9
41767,12
41768,12
41769,15
41770,15
41771,9
41772,12
41773,12
41774,37
41775,9
41776,9
41777,12
41778,47
41779,12
41780,0
41781,12
41782,0
41783,12
41784,12
41785,12
41786,0
41787,12
41788,0
41789,12
41790,47
41791,15
41792,53
41793,53
41794,53
41795,15
41796,53
41797,15
41798,53
41799,15
41800,53
41801,53
41802,53
41803,15
41804,53
41805,15
41806,53
41807,15
41808,15
41809,37
41810,37
41811,47
41812,53
41813,53
41814,37
41815,47
41816,53
41817,53
41818,37
41819,18
41820,18
41821,47
41822,53
41823,53
41824,37
41825,37
41826,47
41827,15
41828,15
41829,12
41830,12
41831,12
41832,12
41833,19
41834,19
41835,19
41836,19
41837,12
41838,12
41839,12
41840,12
41841,12
41842,12
41843,15
41844,53
41845,53
41846,37
41847,12
41848,15
41849,15
41850,12
41851,12
41852,37
41853,53
41854,53
41855,37
41856,19
41857,19
41858,15
41859,15
41860,15
41861,53
41862,53
41863,37
41864,19
41865,19
41866,15
41867,15
41868,15
41869,12
41870,12
41871,12
41872,12
41873,53
41874,14
41875,53
41876,14
41877,37
41878,14
41879,53
41880,53
41881,37
41882,15
41883,15
41884,15
41885,37
41886,37
41887,49
41888,15
41889,15
41890,53
41891,53
41892,15
41893,14
41894,37
41895,14
41896,37
41897,15
41898,15
41899,15
41900,15
41901,15
41902,15
41903,3
41904,3
41905,3
41906,3
41907,3
41908,3
41909,37
41910,37
41911,37
41912,3
41913,3
41914,32
41915,32
41916,32
41917,32
41918,32
41919,54
41920,54
41921,19
41922,32
41923,6
41924,32
41925,6
41926,54
41927,54
41928,19
41929,11
41930,11
41931,19
41932,19
41933,19
41934,19
41935,19
41936,19
41937,49
41938,19
41939,19
41940,19
41941,27
41942,27
41943,37
41944,37
41945,37
41946,32
41947,29
41948,29
41949,32
41950,29
41951,29
41952,32
41953,33
41954,33
41955,54
41956,54
41957,29
41958,29
41959,29
41960,37
41961,37
41962,27
41963,27
41964,27
41965,27
41966,33
41967,33
41968,27
41969,27
41970,15
41971,15
41972,15
41973,15
41974,15
41975,3
41976,3
41977,3
41978,3
41979,3
41980,15
41981,15
41982,18
41983,15
41984,3
41985,3
41986,18
41987,15
41988,15
41989,3
41990,3
41991,3
41992,3
41993,15
41994,15
41995,3
41996,3
41997,18
41998,15
41999,15
42000,18
42001,3
42002,34
42003,34
42004,55
42005,1
42006,55
42007,1
42008,3
42009,33
42010,55
42011,55
42012,37
42013,33
42014,55
42015,55
42016,37
42017,11
42018,55
42019,55
42020,37
42021,11
42022,55
42023,55
42024,37
42025,11
42026,55
42027,55
42028,37
42029,12
42030,12
42031,12
42032,49
42033,49
42034,49
42035,49
42036,6
42037,32
42038,53
42039,53
42040,6
42041,32
42042,53
42043,53
42044,6
42045,32
42046,49
42047,49
42048,49
42049,53
42050,49
42051,53
42052,6
42053,6
42054,6
42055,49
42056,49
42057,49
42058,49
42059,6
42060,19
42061,19
42062,6
42063,6
42064,19
42065,19
42066,19
42067,12
42068,12
42069,15
42070,55
42071,15
42072,55
42073,37
42074,15
42075,15
42076,15
42077,19
42078,55
42079,55
42080,37
42081,55
42082,55
42083,55
42084,55
42085,37
42086,37
42087,37
42088,6
42089,6
42090,55
42091,37
42092,55
42093,55
42094,33
42095,55
42096,55
42097,37
42098,9
42099,12
42100,12
42101,33
42102,55
42103,55
42104,37
42105,37
42106,37
42107,19
42108,19
42109,9
42110,12
42111,12
42112,37
42113,55
42114,55
42115,37
42116,32
42117,55
42118,55
42119,12
42120,32
42121,55
42122,55
42123,12
42124,12
42125,12
42126,12
42127,12
42128,12
42129,12
42130,15
42131,15
42132,12
42133,19
42134,55
42135,55
42136,12
42137,15
42138,15
42139,12
42140,19
42141,19
42142,12
42143,12
42144,12
42145,12
42146,12
42147,12
42148,12
42149,55
42150,55
42151,55
42152,55
42153,55
42154,15
42155,15
42156,55
42157,15
42158,15
42159,15
42160,14
42161,14
42162,14
42163,37
42164,3
42165,3
42166,3
42167,3
42168,3
42169,3
42170,6
42171,6
42172,37
42173,3
42174,3
42175,3
42176,3
42177,3
42178,6
42179,6
42180,55
42181,3
42182,55
42183,3
42184,55
42185,3
42186,3
42187,6
42188,6
42189,55
42190,3
42191,3
42192,55
42193,55
42194,55
42195,37
42196,32
42197,11
42198,11
42199,27
42200,19
42201,11
42202,11
42203,27
42204,27
42205,32
42206,32
42207,27
42208,19
42209,11
42210,11
42211,19
42212,11
42213,11
42214,19
42215,11
42216,11
42217,19
42218,11
42219,6
42220,6
42221,11
42222,27
42223,27
42224,33
42225,33
42226,33
42227,29
42228,29
42229,29
42230,49
42231,29
42232,29
42233,29
42234,27
42235,27
42236,33
42237,33
42238,27
42239,27
42240,33
42241,33
42242,27
42243,33
42244,27
42245,27
42246,47
42247,47
42248,47
42249,47
42250,47
42251,1
42252,15
42253,15
42254,15
42255,15
42256,15
42257,3
42258,18
42259,18
42260,15
42261,15
42262,18
42263,15
42264,18
42265,18
42266,15
42267,15
42268,18
42269,1
42270,1
42271,3
42272,3
42273,55
42274,55
42275,3
42276,55
42277,55
42278,55
42279,37
42280,37
42281,55
42282,55
42283,37
42284,37
42285,55
42286,55
42287,37
42288,32
42289,12
42290,12
42291,39
42292,39
42293,6
42294,12
42295,12
42296,12
42297,12
42298,39
42299,39
42300,32
42301,6
42302,32
42303,32
42304,6
42305,32
42306,53
42307,53
42308,6
42309,32
42310,53
42311,53
42312,6
42313,32
42314,49
42315,49
42316,49
42317,49
42318,6
42319,18
42320,18
42321,19
42322,37
42323,12
42324,12
42325,15
42326,55
42327,15
42328,55
42329,37
42330,55
42331,15
42332,15
42333,19
42334,55
42335,55
42336,37
42337,19
42338,54
42339,54
42340,15
42341,15
42342,37
42343,33
42344,55
42345,55
42346,18
42347,18
42348,55
42349,55
42350,55
42351,55
42352,55
42353,37
42354,37
42355,37
42356,37
42357,37
42358,55
42359,55
42360,55
42361,18
42362,18
42363,9
42364,55
42365,55
42366,33
42367,37
42368,37
42369,37
42370,9
42371,55
42372,55
42373,33
42374,37
42375,37
42376,37
42377,18
42378,18
42379,37
42380,55
42381,55
42382,37
42383,37
42384,55
42385,55
42386,37
42387,9
42388,9
42389,9
42390,55
42391,55
42392,37
42393,9
42394,9
42395,9
42396,49
42397,15
42398,15
42399,37
42400,12
42401,12
42402,12
42403,12
42404,12
42405,12
42406,55
42407,55
42408,37
42409,12
42410,12
42411,12
42412,19
42413,19
42414,55
42415,55
42416,37
42417,37
42418,19
42419,19
42420,12
42421,12
42422,12
42423,19
42424,19
42425,19
42426,55
42427,55
42428,37
42429,55
42430,55
42431,55
42432,55
42433,6
42434,6
42435,6
42436,6
42437,55
42438,55
42439,15
42440,15
42441,55
42442,19
42443,19
42444,15
42445,15
42446,15
42447,15
42448,15
42449,15
42450,37
42451,37
42452,37
42453,6
42454,6
42455,55
42456,3
42457,3
42458,55
42459,3
42460,3
42461,55
42462,3
42463,3
42464,55
42465,3
42466,3
42467,6
42468,6
42469,19
42470,19
42471,55
42472,55
42473,55
42474,37
42475,37
42476,55
42477,37
42478,55
42479,37
42480,37
42481,37
42482,27
42483,32
42484,32
42485,6
42486,6
42487,37
42488,37
42489,32
42490,11
42491,11
42492,27
42493,27
42494,37
42495,19
42496,11
42497,11
42498,19
42499,55
42500,55
42501,37
42502,37
42503,19
42504,11
42505,11
42506,27
42507,27
42508,27
42509,27
42510,33
42511,29
42512,29
42513,33
42514,29
42515,29
42516,33
42517,29
42518,29
42519,49
42520,33
42521,29
42522,29
42523,33
42524,33
42525,33
42526,29
42527,29
42528,54
42529,54
42530,29
42531,49
42532,29
42533,29
42534,54
42535,54
42536,29
42537,33
42538,29
42539,33
42540,29
42541,33
42542,33
42543,54
42544,54
42545,1
42546,1
42547,15
42548,15
42549,1
42550,3
42551,18
42552,18
42553,18
42554,18
42555,18
42556,3
42557,3
42558,3
42559,3
42560,55
42561,55
42562,1
42563,1
42564,3
42565,3
42566,33
42567,33
42568,37
42569,24
42570,12
42571,12
42572,11
42573,11
42574,37
42575,55
42576,55
42577,37
42578,18
42579,18
42580,37
42581,12
42582,11
42583,11
42584,12
42585,12
42586,11
42587,11
42588,37
42589,37
42590,55
42591,55
42592,37
42593,24
42594,32
42595,32
42596,12
42597,32
42598,12
42599,12
42600,12
42601,12
42602,12
42603,32
42604,32
42605,32
42606,12
42607,32
42608,32
42609,32
42610,12
42611,32
42612,12
42613,12
42614,12
42615,48
42616,53
42617,53
42618,12
42619,12
42620,12
42621,12
42622,12
42623,12
42624,12
42625,12
42626,12
42627,18
42628,18
42629,55
42630,12
42631,12
42632,12
42633,12
42634,12
42635,12
42636,12
42637,12
42638,12
42639,55
42640,12
42641,12
42642,55
42643,55
42644,55
42645,55
42646,25
42647,12
42648,55
42649,55
42650,55
42651,55
42652,55
42653,55
42654,12
42655,55
42656,12
42657,55
42658,12
42659,12
42660,55
42661,12
42662,12
42663,19
42664,55
42665,55
42666,55
42667,55
42668,55
42669,55
42670,12
42671,12
42672,37
42673,18
42674,18
42675,37
42676,55
42677,55
42678,37
42679,55
42680,55
42681,37
42682,55
42683,37
42684,55
42685,55
42686,55
42687,37
42688,55
42689,55
42690,55
42691,37
42692,12
42693,12
42694,12
42695,55
42696,55
42697,18
42698,18
42699,37
42700,55
42701,55
42702,55
42703,37
42704,55
42705,55
42706,55
42707,55
42708,55
42709,12
42710,19
42711,55
42712,55
42713,12
42714,12
42715,12
42716,12
42717,12
42718,55
42719,12
42720,12
42721,55
42722,19
42723,12
42724,55
42725,12
42726,55
42727,12
42728,12
42729,12
42730,12
42731,55
42732,55
42733,55
42734,55
42735,55
42736,12
42737,12
42738,55
42739,55
42740,55
42741,55
42742,37
42743,6
42744,6
42745,37
42746,12
42747,12
42748,12
42749,14
42750,55
42751,55
42752,37
42753,19
42754,19
42755,12
42756,55
42757,55
42758,37
42759,6
42760,6
42761,55
42762,3
42763,3
42764,19
42765,19
42766,55
42767,3
42768,3
42769,3
42770,55
42771,3
42772,55
42773,55
42774,3
42775,3
42776,26
42777,19
42778,11
42779,11
42780,26
42781,19
42782,11
42783,11
42784,19
42785,11
42786,11
42787,19
42788,11
42789,11
42790,19
42791,11
42792,11
42793,19
42794,19
42795,37
42796,19
42797,19
42798,19
42799,19
42800,19
42801,19
42802,54
42803,54
42804,19
42805,26
42806,19
42807,19
42808,33
42809,32
42810,32
42811,33
42812,48
42813,33
42814,48
42815,33
42816,27
42817,27
42818,6
42819,6
42820,6
42821,6
42822,6
42823,6
42824,6
42825,6
42826,6
42827,6
42828,6
42829,6
42830,18
42831,18
42832,6
42833,6
42834,18
42835,18
42836,6
42837,18
42838,18
42839,6
42840,18
42841,18
42842,6
42843,6
42844,6
42845,6
42846,6
42847,6
42848,6
42849,6
42850,6
42851,6
42852,1
42853,1
42854,6
42855,6
42856,6
42857,6
42858,29
42859,29
42860,29
42861,29
42862,6
42863,6
42864,29
42865,29
42866,33
42867,33
42868,29
42869,29
42870,15
42871,15
42872,37
42873,37
42874,37
42875,19
42876,49
42877,49
42878,15
42879,15
42880,6
42881,6
42882,6
42883,6
42884,15
42885,6
42886,6
42887,6
42888,6
42889,1
42890,15
42891,15
42892,15
42893,15
42894,15
42895,15
42896,3
42897,3
42898,15
42899,15
42900,18
42901,3
42902,3
42903,3
42904,1
42905,1
42906,3
42907,55
42908,55
42909,55
42910,55
42911,33
42912,12
42913,12
42914,11
42915,11
42916,0
42917,37
42918,11
42919,11
42920,33
42921,55
42922,55
42923,37
42924,33
42925,55
42926,55
42927,37
42928,37
42929,55
42930,55
42931,37
42932,37
42933,37
42934,37
42935,37
42936,55
42937,11
42938,11
42939,37
42940,37
42941,55
42942,55
42943,37
42944,12
42945,12
42946,12
42947,12
42948,32
42949,6
42950,6
42951,32
42952,6
42953,32
42954,32
42955,6
42956,12
42957,12
42958,12
42959,32
42960,32
42961,12
42962,12
42963,6
42964,12
42965,12
42966,12
42967,12
42968,12
42969,12
42970,12
42971,6
42972,32
42973,32
42974,32
42975,6
42976,19
42977,19
42978,55
42979,55
42980,55
42981,12
42982,12
42983,15
42984,15
42985,55
42986,55
42987,55
42988,12
42989,12
42990,15
42991,15
42992,55
42993,55
42994,55
42995,55
42996,55
42997,19
42998,55
42999,55
43000,37
43001,6
43002,6
43003,37
43004,6
43005,6
43006,19
43007,19
43008,9
43009,55
43010,55
43011,32
43012,12
43013,12
43014,37
43015,37
43016,37
43017,32
43018,55
43019,55
43020,37
43021,37
43022,37
43023,37
43024,37
43025,37
43026,37
43027,37
43028,19
43029,19
43030,6
43031,6
43032,6
43033,55
43034,55
43035,55
43036,12
43037,12
43038,14
43039,14
43040,55
43041,6
43042,6
43043,55
43044,55
43045,55
43046,14
43047,14
43048,55
43049,19
43050,19
43051,55
43052,55
43053,55
43054,55
43055,55
43056,55
43057,55
43058,12
43059,12
43060,14
43061,14
43062,55
43063,55
43064,55
43065,55
43066,14
43067,14
43068,55
43069,55
43070,55
43071,55
43072,55
43073,55
43074,55
43075,14
43076,14
43077,55
43078,6
43079,6
43080,55
43081,15
43082,15
43083,37
43084,37
43085,14
43086,37
43087,55
43088,55
43089,37
43090,55
43091,15
43092,15
43093,14
43094,14
43095,14
43096,14
43097,37
43098,19
43099,19
43100,55
43101,15
43102,15
43103,14
43104,14
43105,37
43106,55
43107,15
43108,15
43109,14
43110,14
43111,3
43112,3
43113,55
43114,3
43115,3
43116,6
43117,6
43118,6
43119,6
43120,55
43121,3
43122,3
43123,6
43124,6
43125,6
43126,6
43127,55
43128,37
43129,55
43130,3
43131,3
43132,19
43133,19
43134,55
43135,55
43136,55
43137,32
43138,55
43139,55
43140,32
43141,32
43142,32
43143,32
43144,32
43145,32
43146,32
43147,32
43148,6
43149,6
43150,32
43151,32
43152,32
43153,6
43154,6
43155,55
43156,37
43157,37
43158,37
43159,32
43160,32
43161,32
43162,33
43163,33
43164,33
43165,27
43166,27
43167,1
43168,15
43169,15
43170,15
43171,15
43172,15
43173,1
43174,1
43175,1
43176,1
43177,1
43178,1
43179,3
43180,3
43181,3
43182,3
43183,0
43184,33
43185,33
43186,37
43187,33
43188,33
43189,33
43190,37
43191,37
43192,33
43193,33
43194,33
43195,33
43196,37
43197,12
43198,11
43199,11
43200,12
43201,12
43202,37
43203,37
43204,37
43205,12
43206,11
43207,11
43208,0
43209,0
43210,12
43211,12
43212,12
43213,12
43214,23
43215,37
43216,37
43217,37
43218,37
43219,37
43220,32
43221,32
43222,32
43223,32
43224,32
43225,32
43226,32
43227,32
43228,12
43229,12
43230,12
43231,12
43232,12
43233,15
43234,15
43235,32
43236,32
43237,12
43238,53
43239,53
43240,6
43241,6
43242,32
43243,49
43244,49
43245,49
43246,49
43247,37
43248,19
43249,19
43250,19
43251,37
43252,18
43253,18
43254,37
43255,19
43256,19
43257,19
43258,19
43259,12
43260,12
43261,12
43262,37
43263,37
43264,37
43265,18
43266,18
43267,12
43268,12
43269,12
43270,37
43271,37
43272,37
43273,37
43274,12
43275,12
43276,12
43277,12
43278,12
43279,12
43280,9
43281,12
43282,12
43283,32
43284,32
43285,32
43286,37
43287,32
43288,32
43289,32
43290,37
43291,18
43292,18
43293,37
43294,32
43295,32
43296,37
43297,47
43298,32
43299,32
43300,37
43301,47
43302,9
43303,9
43304,37
43305,9
43306,9
43307,0
43308,0
43309,47
43310,53
43311,53
43312,37
43313,9
43314,9
43315,9
43316,53
43317,53
43318,37
43319,18
43320,18
43321,9
43322,9
43323,9
43324,19
43325,19
43326,32
43327,15
43328,32
43329,15
43330,32
43331,12
43332,19
43333,19
43334,19
43335,19
43336,12
43337,19
43338,19
43339,12
43340,12
43341,56
43342,56
43343,37
43344,14
43345,14
43346,14
43347,37
43348,19
43349,19
43350,19
43351,19
43352,14
43353,14
43354,14
43355,37
43356,37
43357,37
43358,37
43359,18
43360,18
43361,3
43362,3
43363,3
43364,37
43365,18
43366,18
43367,3
43368,3
43369,3
43370,18
43371,18
43372,3
43373,3
43374,3
43375,3
43376,3
43377,3
43378,3
43379,3
43380,3
43381,32
43382,32
43383,32
43384,18
43385,18
43386,37
43387,19
43388,32
43389,32
43390,49
43391,19
43392,32
43393,6
43394,32
43395,6
43396,32
43397,32
43398,19
43399,32
43400,32
43401,54
43402,54
43403,19
43404,32
43405,32
43406,19
43407,19
43408,6
43409,19
43410,6
43411,54
43412,54
43413,19
43414,6
43415,6
43416,54
43417,54
43418,1
43419,1
43420,15
43421,15
43422,1
43423,3
43424,3
43425,15
43426,15
43427,3
43428,49
43429,35
43430,35
43431,35
43432,35
43433,35
43434,35
43435,35
43436,32
43437,49
43438,49
43439,49
43440,49
43441,49
43442,32
43443,46
43444,46
43445,32
43446,32
43447,32
43448,32
43449,49
43450,32
43451,17
43452,17
43453,49
43454,17
43455,17
43456,17
43457,49
43458,17
43459,17
43460,17
43461,17
43462,17
43463,17
43464,17
43465,17
43466,17
43467,17
43468,15
43469,15
43470,17
43471,19
43472,19
43473,17
43474,17
43475,17
43476,17
43477,17
43478,15
43479,15
43480,17
43481,19
43482,19
43483,19
43484,19
43485,17
43486,54
43487,54
43488,17
43489,17
43490,17
43491,17
43492,37
43493,37
43494,19
43495,19
43496,55
43497,55
43498,55
43499,55
43500,55
43501,55
43502,55
43503,55
43504,55
43505,33
43506,49
43507,55
43508,49
43509,55
43510,55
43511,49
43512,55
43513,49
43514,33
43515,9
43516,55
43517,55
43518,33
43519,55
43520,55
43521,37
43522,37
43523,37
43524,9
43525,9
43526,33
43527,55
43528,55
43529,55
43530,55
43531,9
43532,33
43533,55
43534,55
43535,9
43536,33
43537,9
43538,55
43539,55
43540,55
43541,55
43542,9
43543,49
43544,12
43545,12
43546,12
43547,19
43548,19
43549,55
43550,19
43551,19
43552,19
43553,19
43554,55
43555,55
43556,55
43557,19
43558,19
43559,55
43560,14
43561,14
43562,14
43563,55
43564,37
43565,37
43566,19
43567,19
43568,55
43569,6
43570,6
43571,1
43572,1
43573,37
43574,37
43575,6
43576,6
43577,19
43578,19
43579,17
43580,1
43581,1
43582,17
43583,17
43584,17
43585,0
43586,0
43587,17
43588,17
43589,17
43590,14
43591,14
43592,37
43593,37
43594,37
43595,17
43596,17
43597,17
43598,14
43599,14
43600,49
43601,17
43602,35
43603,35
43604,17
43605,35
43606,35
43607,17
43608,35
43609,17
43610,35
43611,17
43612,17
43613,35
43614,35
43615,49
43616,17
43617,35
43618,35
43619,17
43620,35
43621,35
43622,14
43623,14
43624,14
43625,14
43626,14
43627,14
43628,14
43629,37
43630,17
43631,17
43632,17
43633,14
43634,14
43635,33
43636,35
43637,35
43638,33
43639,33
43640,1
43641,1
43642,1
43643,1
43644,1
43645,1
43646,3
43647,3
43648,3
43649,15
43650,15
43651,3
43652,1
43653,17
43654,17
43655,17
43656,17
43657,17
43658,17
43659,17
43660,17
43661,35
43662,35
43663,35
43664,35
43665,35
43666,32
43667,32
43668,32
43669,39
43670,32
43671,32
43672,32
43673,39
43674,17
43675,17
43676,17
43677,54
43678,54
43679,17
43680,17
43681,17
43682,17
43683,17
43684,17
43685,17
43686,17
43687,55
43688,55
43689,55
43690,55
43691,55
43692,55
43693,55
43694,55
43695,37
43696,37
43697,55
43698,55
43699,37
43700,37
43701,55
43702,37
43703,37
43704,55
43705,49
43706,9
43707,9
43708,37
43709,33
43710,55
43711,55
43712,37
43713,19
43714,19
43715,55
43716,14
43717,14
43718,14
43719,55
43720,14
43721,14
43722,14
43723,14
43724,14
43725,14
43726,14
43727,14
43728,37
43729,37
43730,14
43731,37
43732,37
43733,37
43734,1
43735,55
43736,55
43737,1
43738,1
43739,1
43740,1
43741,1
43742,37
43743,37
43744,37
43745,17
43746,17
43747,17
43748,17
43749,17
43750,17
43751,35
43752,35
43753,17
43754,17
43755,17
43756,35
43757,35
43758,55
43759,35
43760,35
43761,35
43762,35
43763,35
43764,35
43765,14
43766,14
43767,49
43768,35
43769,35
43770,35
43771,35
43772,35
43773,35
43774,14
43775,14
43776,1
43777,1
43778,1
43779,1
43780,1
43781,1
43782,17
43783,1
43784,1
43785,17
43786,17
43787,17
43788,17
43789,17
43790,17
43791,17
43792,17
43793,17
43794,17
43795,17
43796,17
43797,17
43798,17
43799,17
43800,1
43801,17
43802,17
43803,17
43804,17
43805,17
43806,1
43807,17
43808,17
43809,17
43810,17
43811,17
43812,17
43813,17
43814,17
43815,17
43816,17
43817,39
43818,17
43819,17
43820,17
43821,17
43822,17
43823,17
43824,17
43825,39
43826,39
43827,17
43828,19
43829,19
43830,17
43831,17
43832,17
43833,17
43834,17
43835,17
43836,17
43837,55
43838,55
43839,55
43840,12
43841,12
43842,1
43843,1
43844,55
43845,33
43846,55
43847,55
43848,55
43849,55
43850,55
43851,55
43852,55
43853,55
43854,55
43855,55
43856,55
43857,55
43858,12
43859,55
43860,12
43861,55
43862,55
43863,55
43864,55
43865,1
43866,1
43867,19
43868,19
43869,55
43870,55
43871,55
43872,55
43873,33
43874,55
43875,55
43876,55
43877,33
43878,12
43879,12
43880,55
43881,33
43882,55
43883,55
43884,55
43885,55
43886,55
43887,55
43888,55
43889,55
43890,55
43891,55
43892,55
43893,55
43894,55
43895,12
43896,19
43897,19
43898,12
43899,55
43900,55
43901,55
43902,55
43903,55
43904,55
43905,14
43906,55
43907,55
43908,55
43909,19
43910,19
43911,19
43912,19
43913,14
43914,14
43915,14
43916,55
43917,55
43918,14
43919,14
43920,6
43921,6
43922,37
43923,17
43924,17
43925,17
43926,1
43927,17
43928,17
43929,17
43930,17
43931,17
43932,17
43933,17
43934,17
43935,17
43936,17
43937,17
43938,39
43939,39
43940,17
43941,17
43942,17
43943,55
43944,17
43945,35
43946,35
43947,19
43948,19
43949,37
43950,17
43951,17
43952,17
43953,17
43954,17
43955,17
43956,14
43957,14
43958,17
43959,17
43960,17
43961,14
43962,14
43963,26
43964,35
43965,33
43966,33
43967,35
43968,35
43969,33
43970,35
43971,35
43972,14
43973,14
43974,35
43975,33
43976,35
43977,35
43978,33
43979,33
43980,3
43981,3
43982,3
43983,15
43984,15
43985,3
43986,17
43987,1
43988,1
43989,17
43990,17
43991,17
43992,1
43993,1
43994,1
43995,1
43996,1
43997,17
43998,17
43999,17
44000,17
44001,17
44002,17
44003,17
44004,55
44005,35
44006,35
44007,35
44008,35
44009,35
44010,35
44011,35
44012,37
44013,35
44014,37
44015,35
44016,35
44017,35
44018,35
44019,32
44020,39
44021,39
44022,35
44023,32
44024,49
44025,49
44026,35
44027,35
44028,35
44029,35
44030,19
44031,19
44032,17
44033,17
44034,17
44035,17
44036,17
44037,17
44038,17
44039,17
44040,17
44041,17
44042,37
44043,37
44044,55
44045,55
44046,55
44047,55
44048,55
44049,9
44050,9
44051,35
44052,55
44053,35
44054,35
44055,35
44056,55
44057,55
44058,9
44059,9
44060,35
44061,35
44062,9
44063,35
44064,35
44065,55
44066,55
44067,55
44068,32
44069,55
44070,55
44071,55
44072,6
44073,6
44074,55
44075,55
44076,55
44077,55
44078,55
44079,55
44080,55
44081,55
44082,14
44083,55
44084,55
44085,55
44086,14
44087,14
44088,14
44089,55
44090,55
44091,14
44092,14
44093,14
44094,55
44095,14
44096,14
44097,55
44098,55
44099,14
44100,55
44101,55
44102,55
44103,35
44104,35
44105,55
44106,35
44107,35
44108,35
44109,35
44110,55
44111,35
44112,35
44113,55
44114,35
44115,35
44116,35
44117,35
44118,55
44119,35
44120,35
44121,55
44122,55
44123,55
44124,35
44125,35
44126,35
44127,35
44128,35
44129,35
44130,35
44131,35
44132,55
44133,1
44134,17
44135,17
44136,17
44137,17
44138,17
44139,1
44140,1
44141,1
44142,12
44143,12
44144,37
44145,37
44146,37
44147,33
44148,33
44149,33
44150,37
44151,12
44152,33
44153,33
44154,12
44155,12
44156,37
44157,37
44158,37
44159,9
44160,12
44161,12
44162,12
44163,12
44164,37
44165,37
44166,37
44167,49
44168,49
44169,49
44170,1
44171,1
44172,37
44173,14
44174,14
44175,14
44176,14
44177,14
44178,14
44179,12
44180,12
44181,12
44182,14
44183,14
44184,14
44185,14
44186,14
44187,17
44188,1
44189,1
44190,1
44191,1
44192,1
44193,1
44194,17
44195,17
44196,17
44197,14
44198,14
44199,14
44200,14
44201,14
44202,14
44203,14
44204,14
44205,49
44206,49
44207,17
44208,17
44209,17
44210,14
44211,14
44212,14
44213,14
44214,14
44215,14
44216,14
44217,14
44218,14
44219,55
44220,55
44221,55
44222,55
44223,14
44224,14
44225,17
44226,1
44227,1
44228,14
44229,14
44230,37
44231,35
44232,35
44233,35
44234,14
44235,14
44236,35
44237,35
44238,35
44239,35
44240,35
44241,35
44242,55
44243,12
44244,12
44245,37
44246,37
44247,55
44248,9
44249,35
44250,35
44251,35
44252,35
44253,55
44254,12
44255,12
44256,12
44257,12
44258,33
44259,33
44260,33
44261,14
44262,14
44263,33
44264,33
44265,33
44266,33
44267,33
44268,33
44269,1
44270,1
44271,1
44272,1
44273,1
44274,1
44275,14
44276,14
44277,14
44278,14
44279,14
44280,35
44281,35
44282,1
44283,1
44284,1
44285,1
44286,1
44287,1
44288,55
44289,55
44290,55
44291,1
44292,1
44293,55
44294,17
44295,1
44296,1
44297,14
44298,14
44299,14
44300,14
44301,14
44302,14
44303,14
44304,14
44305,17
44306,35
44307,35
44308,14
44309,14
44310,35
44311,35
44312,35
44313,35
44314,35
44315,35
44316,35
44317,35
44318,35
44319,35
44320,35
44321,17
44322,39
44323,39
44324,39
44325,39
44326,17
44327,17
44328,17
44329,17
44330,17
44331,17
44332,55
44333,37
44334,37
44335,55
44336,55
44337,55
44338,55
44339,12
44340,12
44341,37
44342,37
44343,55
44344,55
44345,55
44346,55
44347,12
44348,12
44349,14
44350,55
44351,55
44352,55
44353,55
44354,55
44355,55
44356,14
44357,14
44358,14
44359,14
44360,55
44361,55
44362,55
44363,55
44364,14
44365,14
44366,24
44367,14
44368,14
44369,14
44370,14
44371,14
44372,14
44373,14
44374,14
44375,14
44376,14
44377,24
44378,17
44379,14
44380,14
44381,14
44382,14
44383,55
44384,17
44385,17
44386,17
44387,14
44388,14
44389,14
44390,14
44391,14
44392,35
44393,35
44394,35
44395,14
44396,14
44397,14
44398,14
44399,33
44400,33
44401,33
44402,35
44403,35
44404,35
44405,14
44406,14
44407,29
44408,14
44409,14
44410,14
44411,14
44412,6
44413,1
44414,35
44415,35
44416,14
44417,14
44418,19
44419,6
44420,6
44421,15
44422,15
44423,6
44424,6
44425,37
44426,37
44427,6
44428,6
44429,19
44430,49
44431,49
44432,49
44433,49
44434,37
44435,19
44436,35
44437,49
44438,49
44439,35
44440,35
44441,49
44442,49
44443,37
44444,46
44445,6
44446,6
44447,49
44448,49
44449,15
44450,15
44451,3
44452,3
44453,3
44454,3
44455,32
44456,55
44457,55
44458,55
44459,55
44460,35
44461,35
44462,35
44463,35
44464,55
44465,55
44466,55
44467,55
44468,35
44469,35
44470,35
44471,35
44472,55
44473,35
44474,35
44475,35
44476,35
44477,55
44478,35
44479,35
44480,35
44481,35
44482,35
44483,17
44484,17
44485,17
44486,1
44487,1
44488,17
44489,17
44490,17
44491,17
44492,17
44493,17
44494,17
44495,17
44496,17
44497,17
44498,17
44499,17
44500,17
44501,17
44502,17
44503,1
44504,1
44505,1
44506,33
44507,37
44508,37
44509,9
44510,12
44511,12
44512,12
44513,12
44514,14
44515,14
44516,14
44517,14
44518,14
44519,35
44520,35
44521,35
44522,35
44523,35
44524,35
44525,35
44526,35
44527,35
44528,35
44529,35
44530,35
44531,35
44532,35
44533,35
44534,35
44535,35
44536,35
44537,35
44538,17
44539,39
44540,39
44541,39
44542,39
44543,17
44544,0
44545,0
44546,0
44547,14
44548,14
44549,37
44550,17
44551,17
44552,17
44553,14
44554,14
44555,17
44556,17
44557,17
44558,14
44559,14
44560,3
44561,3
44562,3
44563,15
44564,15
44565,3
44566,32
44567,12
44568,12
44569,55
44570,55
44571,55
44572,19
44573,19
44574,14
44575,14
44576,14
44577,14
44578,14
44579,14
44580,17
44581,17
44582,17
44583,55
44584,55
44585,37
44586,14
44587,14
44588,14
44589,32
44590,32
44591,14
44592,19
44593,19
44594,14
44595,37
44596,37
44597,32
44598,33
44599,35
44600,35
44601,33
44602,33
44603,35
44604,33
44605,33
44606,35
44607,35
44608,35
44609,35
44610,35
44611,35
44612,35
44613,35
44614,35
44615,35
44616,35
44617,35
44618,35
44619,35
44620,17
44621,17
44622,17
44623,39
44624,39
44625,17
44626,17
44627,17
44628,17
44629,17
44630,17
44631,55
44632,1
44633,1
44634,12
44635,12
44636,14
44637,14
44638,17
44639,17
44640,17
44641,14
44642,14
